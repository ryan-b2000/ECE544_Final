
`timescale 1 ps / 1 ps

module n4fpga
(
   input				clk,				// 100Mhz clock input
   input                btnC,            	// center pushbutton
   input                btnU,            	// UP (North) pusbhbutton
   input                btnL,            	// LEFT (West) pushbutton
   input                btnD,           	// DOWN (South) pushbutton  - used for system reset
   input                btnR,            	// RIGHT (East) pushbutton
   input                btnCpuReset,    	// CPU reset pushbutton
   input    [15:0]      sw,                 // slide switches on Nexys 4
   output   [15:0]     led,            	// LEDs on Nexys 4  
   
   
   output [7:0]        an,             		// Seven Segment display
   output [6:0]        seg,					// Digits
   output              dp,             		// decimal point display on the seven segment 
   
   input                uart_rtl_rxd,    // USB UART Rx and Tx on Nexys 4
   output               uart_rtl_txd,     
    
   inout     [7:0]       JA,             // JA PmodOLED connector 
  // inout     [2:0]       JC,             // JC PMODHB3 connector
  // inout    [7:0]        JD,             // JD PmodENC connector
   
   //Pin assignments of the DDR3 Module generated by MIG7 IP
   output [12:0] ddr2_sdram_addr,       
   output [2:0]ddr2_sdram_ba,
   output ddr2_sdram_cas_n,
   output [0:0]ddr2_sdram_ck_n,
   output [0:0]ddr2_sdram_ck_p,
   output [0:0]ddr2_sdram_cke,
   output [0:0]ddr2_sdram_cs_n,
   output [1:0]ddr2_sdram_dm,
   inout [15:0]ddr2_sdram_dq,
   inout [1:0]ddr2_sdram_dqs_n,
   inout [1:0]ddr2_sdram_dqs_p,
   output [0:0]ddr2_sdram_odt,
   output ddr2_sdram_ras_n,
   output ddr2_sdram_we_n
  );


// internal variables
// System Clock and Reset 
logic   sysclk;            
logic   sysreset_n, sysreset;
logic   sys_clock;
logic   reset;



wire [15:0]DDR2_0_dq;
wire [12:0]DDR2_0_addr;
wire [2:0]DDR2_0_ba;
wire [1:0]DDR2_0_dm;
wire [1:0]DDR2_0_dqs_n;
wire [1:0]DDR2_0_dqs_p;

wire DDR2_0_cas_n, DDR2_0_ck_n, DDR2_0_ck_p, DDR2_0_cke, DDR2_0_cs_n, DDR2_0_odt, DDR2_0_ras_n, DDR2_0_we_n;

wire [15:0]GPIO_0_IN_tri_i;
wire [15:0]GPIO_0_OUT_tri_o;

wire SPI_io0_i, SPI_io0_io, SPI_io0_o, SPI_io0_t;
wire SPI_io1_i, SPI_io1_io, SPI_io1_o, SPI_io1_t;
wire SPI_sck_i, SPI_sck_io, SPI_sck_o, SPI_sck_t;
wire SPI_ss_i, SPI_ss_io, SPI_ss_o, SPI_ss_t;

wire UART_0_rxd, UART_0_txd;




// SPI Interface
//logic acl_spi_io0_i, acl_spi_io0_io, acl_spi_io0_o, acl_spi_io0_t;
//logic acl_spi_io1_i, acl_spi_io1_io, acl_spi_io1_o, acl_spi_io1_t;
//logic acl_spi_sck_i, acl_spi_sck_io, acl_spi_sck_o, acl_spi_sck_t;
//logic acl_spi_ss_i,  acl_spi_ss_io,  acl_spi_ss_o,  acl_spi_ss_t;

// DIP Switches
//logic [15:0]dip_switches_tri_i;

// Switch LED GPIOs
//logic switch_leds_tri_i_0, switch_leds_tri_io_0, switch_leds_tri_o_0, switch_leds_tri_t_0;
//logic switch_leds_tri_i_1, switch_leds_tri_io_1, switch_leds_tri_o_1, switch_leds_tri_t_1; 
//logic switch_leds_tri_i_2, switch_leds_tri_io_2, switch_leds_tri_o_2, switch_leds_tri_t_2; 
//logic switch_leds_tri_i_3, switch_leds_tri_io_3, switch_leds_tri_o_3, switch_leds_tri_t_3; 
//logic switch_leds_tri_i_4, switch_leds_tri_io_4, switch_leds_tri_o_4, switch_leds_tri_t_4; 
//logic switch_leds_tri_i_5, switch_leds_tri_io_5, switch_leds_tri_o_5, switch_leds_tri_t_5; 
//logic switch_leds_tri_i_6, switch_leds_tri_io_6, switch_leds_tri_o_6, switch_leds_tri_t_6; 
//logic switch_leds_tri_i_7, switch_leds_tri_io_7, switch_leds_tri_o_7, switch_leds_tri_t_7; 
//logic switch_leds_tri_i_8, switch_leds_tri_io_8, switch_leds_tri_o_8, switch_leds_tri_t_8; 
//logic switch_leds_tri_i_9, switch_leds_tri_io_9, switch_leds_tri_o_9, switch_leds_tri_t_9; 
//logic switch_leds_tri_i_10, switch_leds_tri_io_10, switch_leds_tri_o_10, switch_leds_tri_t_10; 
//logic switch_leds_tri_i_11, switch_leds_tri_io_11, switch_leds_tri_o_11, switch_leds_tri_t_11; 
//logic switch_leds_tri_i_12, switch_leds_tri_io_12, switch_leds_tri_o_12, switch_leds_tri_t_12; 
//logic switch_leds_tri_i_13, switch_leds_tri_io_13, switch_leds_tri_o_13, switch_leds_tri_t_13; 
//logic switch_leds_tri_i_14, switch_leds_tri_io_14, switch_leds_tri_o_14, switch_leds_tri_t_14;
//logic switch_leds_tri_i_15, switch_leds_tri_io_15, switch_leds_tri_o_15, switch_leds_tri_t_15;

// Rotary encoder pins
//logic 	Pmod_out_0_pin1_i, Pmod_out_0_pin1_io, Pmod_out_0_pin1_o, Pmod_out_0_pin1_t;
//logic 	Pmod_out_0_pin2_i, Pmod_out_0_pin2_io, Pmod_out_0_pin2_o, Pmod_out_0_pin2_t;
//logic 	Pmod_out_0_pin3_i, Pmod_out_0_pin3_io, Pmod_out_0_pin3_o, Pmod_out_0_pin3_t;
//logic 	Pmod_out_0_pin4_i, Pmod_out_0_pin4_io, Pmod_out_0_pin4_o, Pmod_out_0_pin4_t;
//logic 	Pmod_out_0_pin7_i, Pmod_out_0_pin7_io, Pmod_out_0_pin7_o, Pmod_out_0_pin7_t; 
//logic 	Pmod_out_0_pin8_i, Pmod_out_0_pin8_io, Pmod_out_0_pin8_o, Pmod_out_0_pin8_t; 
//logic 	Pmod_out_0_pin9_i, Pmod_out_0_pin9_io, Pmod_out_0_pin9_o, Pmod_out_0_pin9_t;
//logic 	Pmod_out_0_pin10_i,Pmod_out_0_pin10_io, Pmod_out_0_pin10_o, Pmod_out_0_pin10_t;

// OLED pins 
//logic 	PmodOLEDrgb_out_0_pin1_i, PmodOLEDrgb_out_0_pin1_io, PmodOLEDrgb_out_0_pin1_o, PmodOLEDrgb_out_0_pin1_t; 
//logic 	PmodOLEDrgb_out_0_pin2_i, PmodOLEDrgb_out_0_pin2_io, PmodOLEDrgb_out_0_pin2_o, PmodOLEDrgb_out_0_pin2_t; 
//logic 	PmodOLEDrgb_out_0_pin3_i, PmodOLEDrgb_out_0_pin3_io, PmodOLEDrgb_out_0_pin3_o, PmodOLEDrgb_out_0_pin3_t; 
//logic 	PmodOLEDrgb_out_0_pin4_i, PmodOLEDrgb_out_0_pin4_io, PmodOLEDrgb_out_0_pin4_o, PmodOLEDrgb_out_0_pin4_t; 
//logic 	PmodOLEDrgb_out_0_pin7_i, PmodOLEDrgb_out_0_pin7_io, PmodOLEDrgb_out_0_pin7_o, PmodOLEDrgb_out_0_pin7_t; 
//logic 	PmodOLEDrgb_out_0_pin8_i, PmodOLEDrgb_out_0_pin8_io, PmodOLEDrgb_out_0_pin8_o, PmodOLEDrgb_out_0_pin8_t; 
//logic 	PmodOLEDrgb_out_0_pin9_i, PmodOLEDrgb_out_0_pin9_io, PmodOLEDrgb_out_0_pin9_o, PmodOLEDrgb_out_0_pin9_t; 
//logic 	PmodOLEDrgb_out_0_pin10_i, PmodOLEDrgb_out_0_pin10_io, PmodOLEDrgb_out_0_pin10_o, PmodOLEDrgb_out_0_pin10_t;



// system-wide signals
assign sysclk = clk;
assign sysreset_n = btnCpuReset;        // The CPU reset pushbutton is asserted low.  The other pushbuttons are asserted high
                                      // but the Microblaze for Nexys 4 expects reset to be asserted low
assign sysreset = ~sysreset_n;          // Generate a reset signal that is asserted high for any logic blocks expecting it.

//Debounce module instatiation to control the push button 
//debounce debounce(sysclk,{btnC,btnD,btnU,btnL,btnR},sw,{btnC_W,btnD_W,btnU_W,btnL_W,btnR_W},switch);


assign JA[0] = SPI_io0_io;
assign JA[1] = SPI_io1_io;
assign JA[2] = SPI_sck_io;
assign JA[3] = SPI_ss_io;


// Pmod OLED connections 
//assign JA[0] = PmodOLEDrgb_out_0_pin1_io;
//assign JA[1] = PmodOLEDrgb_out_0_pin2_io;
//assign JA[2] = PmodOLEDrgb_out_0_pin3_io;
//assign JA[3] = PmodOLEDrgb_out_0_pin4_io;
//assign JA[4] = PmodOLEDrgb_out_0_pin7_io;
//assign JA[5] = PmodOLEDrgb_out_0_pin8_io;
//assign JA[6] = PmodOLEDrgb_out_0_pin9_io;
//assign JA[7] = PmodOLEDrgb_out_0_pin10_io;

//assign sw = dip_switches_tri_i;

//assign led[3:0] = {switch_leds_tri_io_3, switch_leds_tri_io_2, switch_leds_tri_io_1, switch_leds_tri_io_0};
//assign led[7:4] = {switch_leds_tri_io_7, switch_leds_tri_io_6, switch_leds_tri_io_5, switch_leds_tri_io_4};
//assign led[11:8] = {switch_leds_tri_io_11, switch_leds_tri_io_10, switch_leds_tri_io_9, switch_leds_tri_io_8};
//assign led[15:12] = {switch_leds_tri_io_15, switch_leds_tri_io_14, switch_leds_tri_io_13, switch_leds_tri_io_12};

// PmodENC signals
// JD - top row
// Pins are assigned such that turning the knob to the right
// causes the rotary count to increment.

embsys embsys_i
   (
    // System Clock and Reset
    .sysclk(sysclk),
    .sysreset(sysreset),
    // DDR2 Signals
    .DDR2_0_addr(ddr2_sdram_addr),
    .DDR2_0_ba(ddr2_sdram_ba),
    .DDR2_0_cas_n(ddr2_sdram_cas_n),
    .DDR2_0_ck_n(ddr2_sdram_ck_n),
    .DDR2_0_ck_p(ddr2_sdram_ck_p),
    .DDR2_0_cke(ddr2_sdram_cke),
    .DDR2_0_cs_n(ddr2_sdram_cs_n),
    .DDR2_0_dm(ddr2_sdram_dm),
    .DDR2_0_dq(ddr2_sdram_dq),
    .DDR2_0_dqs_n(ddr2_sdram_dqs_n),
    .DDR2_0_dqs_p(ddr2_sdram_dqs_p),
    .DDR2_0_odt(ddr2_sdram_odt),
    .DDR2_0_ras_n(ddr2_sdram_ras_n),
    .DDR2_0_we_n(ddr2_sdram_we_n),
    
    .GPIO_0_IN_tri_i(GPIO_0_IN_tri_i),
    .GPIO_0_OUT_tri_o(GPIO_0_OUT_tri_o),
    
    .SPI_io0_i(SPI_io0_i),
    .SPI_io0_o(SPI_io0_o),
    .SPI_io0_t(SPI_io0_t),
    .SPI_io1_i(SPI_io1_i),
    .SPI_io1_o(SPI_io1_o),
    .SPI_io1_t(SPI_io1_t),
    .SPI_sck_i(SPI_sck_i),
    .SPI_sck_o(SPI_sck_o),
    .SPI_sck_t(SPI_sck_t),
    .SPI_ss_i(SPI_ss_i),
    .SPI_ss_o(SPI_ss_o),
    .SPI_ss_t(SPI_ss_t),
    
    .UART_0_rxd(uart_rtl_rxd),
    .UART_0_txd(uart_rtl_txd),
    
    .an_0(an),
    .dp_0(dp),
    .seg_0(seg),
    
    .btnC_0(btnC),
    .btnD_0(btnD),
    .btnL_0(btnL),
    .btnR_0(btnR),
    .btnU_0(btnU),
    
    .led_0(led),
    .sw_0(sw));
        
    
IOBUF SPI_io0_iobuf
     (.I(SPI_io0_o),
      .IO(SPI_io0_io),
      .O(SPI_io0_i),
      .T(SPI_io0_t));
IOBUF SPI_io1_iobuf
     (.I(SPI_io1_o),
      .IO(SPI_io1_io),
      .O(SPI_io1_i),
      .T(SPI_io1_t));
IOBUF SPI_sck_iobuf
     (.I(SPI_sck_o),
      .IO(SPI_sck_io),
      .O(SPI_sck_i),
      .T(SPI_sck_t));
IOBUF SPI_ss_iobuf
     (.I(SPI_ss_o),
      .IO(SPI_ss_io),
      .O(SPI_ss_i),
      .T(SPI_ss_t));
endmodule
